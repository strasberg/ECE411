	mem(0) := To_stdlogicvector(X"02");
	mem(1) := To_stdlogicvector(X"E4");
	mem(2) := To_stdlogicvector(X"80");
	mem(3) := To_stdlogicvector(X"40");
	mem(4) := To_stdlogicvector(X"FF");
	mem(5) := To_stdlogicvector(X"0F");
	mem(6) := To_stdlogicvector(X"61");
	mem(7) := To_stdlogicvector(X"12");
	mem(8) := To_stdlogicvector(X"C0");
	mem(9) := To_stdlogicvector(X"C1");
