--
-- VHDL Architecture ece411.JSRMux.untitled
--
-- Created:
--          by - strasbe1.ews (gelib-057-16.ews.illinois.edu)
--          at - 13:22:41 02/02/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY JSRMux IS
   PORT( 
      clk  : IN     std_logic;
      dest : IN     LC3b_reg;
      sig0 : OUT    std_logic
   );

-- Declarations

END JSRMux ;

--
ARCHITECTURE untitled OF JSRMux IS
BEGIN
END ARCHITECTURE untitled;

